module MM(clk, rst, A, B, N, len, Z);
input clk, rst;
input [31:0] A, B, N;
input [7:0] len;
output [31:0] Z;



endmodule 
