module RL_binary(base, exp, N, R);
input [31:0] base, exp, N;
output [31:0] R;



endmodule
