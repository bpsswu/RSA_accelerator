library verilog;
use verilog.vl_types.all;
entity IO_tb is
end IO_tb;
